package my_uvm_pkg;
    import uvm_pkg::*;
//   `include "driver_interface.sv"
//   `include "monitor_interface.sv"
   `include "packet.sv"
   `include "packet_sequence.sv"
   `include "packet_sequencer.sv"
   `include "packet_driver.sv"
   `include "packet_monitor.sv"
   `include "packet_agent.sv"
   `include "packet_scoreboard.sv"
   `include "packet_env.sv"
   `include "test.sv"
endpackage